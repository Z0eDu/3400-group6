module Grid (
	PIXEL_X,
	PIXEL_Y,
	OUTPUT
);

input  [9:0] PIXEL_X;
input  [9:0] PIXEL_Y;
output [1:0] OUTPUT;

always @(*) begin
	if (PIXEL_X < 

end
